////////////////////////////////////////////////////////////////////////////////
#IGNORE#
#IGNORE#
#IGNORE#
#IGNORE#
////////////////////////////////////////////////////////////////////////////////

module top_const_assign_reversed();
wire [3:0] sink_bus;

assign sink_bus = 4'b0101;
endmodule //top_const_assign_reversed
