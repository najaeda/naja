/* 
  Copyright The Naja Authors.
  SPDX-FileCopyrightText: 2023 The Naja authors <https://github.com/xtofalex/naja/blob/main/AUTHORS>
  SPDX-License-Identifier: Apache-2.0

  Error: referencing bit slice on scalar net.
*/

module model(error, error);
  input error;
  input error;
endmodule

module test();
  model inst(.error(), .error());
endmodule