module model();
endmodule //model

(* PRAGMA1=value1 *)
(* PRAGMA2=value2 *)
(* PRAGMA2 *)
module top(input term);
(* NPRAGMA1=value1 *)
(* NPRAGMA2=value2 *)
(* NPRAGMA2 *)
wire net;

(* IPRAGMA1=value1 *)
(* IPRAGMA2=value2 *)
(* IPRAGMA2 *)
model ins (
);
endmodule //top
