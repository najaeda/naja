module \#model0 (input \%t0 , input \12t1@ , input [3:0] \3 4 , input [-5:2] \## );
endmodule //#model0

module \design@ ();
wire \^n0^ ;
wire \[n1] ;
wire [3:0] \3 4 ;
wire [-5:2] \## ;

\#model0  \0ins  (
  .%t0(\^n0^ ),
  .12t1@(\[n1] ),
  .3 4(\3 4 ),
  .##(\## )
);
endmodule //design@
