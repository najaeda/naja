/*
  Error when instance model does not exist
*/

module test(input i, output o, inout io);
  unknown inst();
endmodule