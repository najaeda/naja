module module2(input a, output c);
endmodule