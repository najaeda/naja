module module1(input a, input b, output c);
endmodule