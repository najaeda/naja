////////////////////////////////////////////////////////////////////////////////
#IGNORE#
#IGNORE#
#IGNORE#
#IGNORE#
////////////////////////////////////////////////////////////////////////////////

module top(input i0, input [31:0] i1, output o, input [31:0] i2, output o_0, output o_1,
 output o_2, output o_3, output o_4, output o_5, output o_6, output o_7, output o_8,
 output o_9, output o_10, output o_11, output o_12, output o_13, output o_14, output o_15,
 output o_16, output o_17, output o_18, output o_19, output o_20, output o_21, output o_22,
 output o_23, output o_24, output o_25, output o_26, output o_27, output o_28, output o_29,
 output o_30, output o_31, output o_32, output o_33, output o_34, output o_35, output o_36,
 output o_37, output o_38, output o_39, output o_40, output o_41, output o_42, output o_43,
 output o_44, output o_45, output o_46, output o_47, output o_48, output o_49, output o_50,
 output o_51, output o_52, output o_53, output o_54, output o_55, output o_56, output o_57,
 output o_58, output o_59, output o_60, output o_61, output o_62, output o_63, output o_64,
 output o_65, output o_66, output o_67, output o_68, output o_69, output o_70, output o_71,
 output o_72, output o_73, output o_74, output o_75, output o_76, output o_77, output o_78,
 output o_79, output o_80, output o_81, output o_82, output o_83, output o_84, output o_85,
 output o_86, output o_87, output o_88, output o_89, output o_90, output o_91, output o_92,
 output o_93, output o_94, output o_95, output o_96, output o_97, output o_98, output o_99,
 output o_100, output o_101, output o_102, output o_103, output o_104, output o_105,
 output o_106, output o_107, output o_108, output o_109, output o_110, output o_111,
 output o_112, output o_113, output o_114, output o_115, output o_116, output o_117,
 output o_118, output o_119, output o_120, output o_121, output o_122, output o_123,
 output o_124, output o_125, output o_126, output o_127, output o_128, output o_129,
 output o_130, output o_131, output o_132, output o_133, output o_134, output o_135,
 output o_136, output o_137, output o_138, output o_139, output o_140, output o_141,
 output o_142, output o_143, output o_144, output o_145, output o_146, output o_147,
 output o_148, output o_149, output o_150, output o_151, output o_152, output o_153,
 output o_154, output o_155, output o_156, output o_157, output o_158, output o_159,
 output o_160, output o_161, output o_162, output o_163, output o_164, output o_165,
 output o_166, output o_167, output o_168, output o_169, output o_170, output o_171,
 output o_172, output o_173, output o_174, output o_175, output o_176, output o_177,
 output o_178, output o_179, output o_180, output o_181, output o_182, output o_183,
 output o_184, output o_185, output o_186, output o_187, output o_188, output o_189,
 output o_190, output o_191, output o_192, output o_193, output o_194, output o_195,
 output o_196, output o_197, output o_198, output o_199);
endmodule //top
