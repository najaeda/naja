////////////////////////////////////////////////////////////////////////////////
#IGNORE#
#IGNORE#
#IGNORE#
#IGNORE#
////////////////////////////////////////////////////////////////////////////////

module AND(input I0, input I1, output Q);
endmodule //AND
module RAM(input CLK, input [31:0] A0, input [31:0] A1, output [127:0] Q);
parameter INVERTED_CLK = "FALSE" ;
parameter WIDTH = 56 ;

endmodule //RAM
