module model();
endmodule //model

(* PRAGMA1="=value1" *)
(* PRAGMA2=12 *)
(* PRAGMA2 *)
module top(input term);
(* NPRAGMA1="=value1" *)
(* NPRAGMA2=88 *)
(* NPRAGMA2 *)
wire net;

(* IPRAGMA1="=value1" *)
(* IPRAGMA2=9 *)
(* IPRAGMA2 *)
model ins (
);
endmodule //top
