////////////////////////////////////////////////////////////////////////////////
#IGNORE#
#IGNORE#
#IGNORE#
#IGNORE#
////////////////////////////////////////////////////////////////////////////////

module top_bus_assign_reversed();
wire [3:0] source_bus;
wire [3:0] sink_bus;

assign sink_bus = source_bus[0:3];
endmodule //top_bus_assign_reversed
