/*
* This is a test file for the auto blackbox generation.
* It contains various test cases to ensure the functionality
* of the blackbox generation process.
*/

module test2();
  wire net0;
  
  auto_blackbox0 ins0(
    .A(net0)
  );

endmodule