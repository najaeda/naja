/*
* This is a test file to test the different conflicting name modules parsin
* policies.
*/

module clash(input A);
  Foo foo();
endmodule

module clash(input B);
endmodule

module Foo();
endmodule

module clash(input C);
endmodule

module clash(input D);
  Foo foo();
endmodule