module top_terms_same_nets(input term0, output [31:0] term1, input [1:1] term2);
endmodule //top_terms_same_nets
