/*
  Error: wire collision
*/

module test();
  wire n0;
  wire n0;
endmodule