////////////////////////////////////////////////////////////////////////////////
#IGNORE#
#IGNORE#
#IGNORE#
#IGNORE#
////////////////////////////////////////////////////////////////////////////////

module top_const_assign_non_contiguous();
wire [5:0] sink_bus;

assign sink_bus[5:4] = 2'b10;

assign sink_bus[2:0] = 3'b101;
endmodule //top_const_assign_non_contiguous
