////////////////////////////////////////////////////////////////////////////////
#IGNORE#
#IGNORE#
#IGNORE#
#IGNORE#
////////////////////////////////////////////////////////////////////////////////

module top(input in, output out);
wire feedtru;

assign feedtru = in;
assign out = feedtru;

endmodule //top
