// SPDX-FileCopyrightText: 2026 The Naja authors <https://github.com/najaeda/naja/blob/main/AUTHORS>
//
// SPDX-License-Identifier: Apache-2.0

module port_directions_top(
  input logic i,
  output logic o,
  inout wire io
);
  assign o = i;
endmodule
