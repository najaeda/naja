////////////////////////////////////////////////////////////////////////////////
#IGNORE#
#IGNORE#
#IGNORE#
#IGNORE#
////////////////////////////////////////////////////////////////////////////////

module top_scalar_assign_output();
wire [1:0] source_bus;
wire scalar_sink;

assign scalar_sink = source_bus[0];
endmodule //top_scalar_assign_output
