module implicit_net0(
    input a,
    input b,
    output y
);
    and and0 (y, a, b, c);
endmodule