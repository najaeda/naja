/*
  Error: referencing bit slice on scalar net.
*/

module model(error, error);
  input error;
  input error;
endmodule

module test();
  model inst(.error(), .error());
endmodule