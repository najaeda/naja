module top();
parameter PARAM0 = 8 ;
parameter PARAM1 = 14 ;

endmodule //top
