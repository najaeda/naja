/*
  Error: unsupported type in instance connection
*/

module test();
  assign n1 = "FOO";
endmodule