/*
  large_hier_gates: synthetic hierarchical gate-level netlist.
*/

module Leaf(input a, input b, input c, output y);
  wire w1, w2, w3, w4;
  and g0(w1, a, b);
  xor g1(w2, w1, c);
  not g2(w3, w2);
  or  g3(w4, w1, w3);
  buf g4(y, w4);
endmodule

module Mid(input [255:0] a, input [255:0] b, input [255:0] c, output [255:0] y);
  Leaf l0(.a(a[0]), .b(b[0]), .c(c[0]), .y(y[0]));
  Leaf l1(.a(a[1]), .b(b[1]), .c(c[1]), .y(y[1]));
  Leaf l2(.a(a[2]), .b(b[2]), .c(c[2]), .y(y[2]));
  Leaf l3(.a(a[3]), .b(b[3]), .c(c[3]), .y(y[3]));
  Leaf l4(.a(a[4]), .b(b[4]), .c(c[4]), .y(y[4]));
  Leaf l5(.a(a[5]), .b(b[5]), .c(c[5]), .y(y[5]));
  Leaf l6(.a(a[6]), .b(b[6]), .c(c[6]), .y(y[6]));
  Leaf l7(.a(a[7]), .b(b[7]), .c(c[7]), .y(y[7]));
  Leaf l8(.a(a[8]), .b(b[8]), .c(c[8]), .y(y[8]));
  Leaf l9(.a(a[9]), .b(b[9]), .c(c[9]), .y(y[9]));
  Leaf l10(.a(a[10]), .b(b[10]), .c(c[10]), .y(y[10]));
  Leaf l11(.a(a[11]), .b(b[11]), .c(c[11]), .y(y[11]));
  Leaf l12(.a(a[12]), .b(b[12]), .c(c[12]), .y(y[12]));
  Leaf l13(.a(a[13]), .b(b[13]), .c(c[13]), .y(y[13]));
  Leaf l14(.a(a[14]), .b(b[14]), .c(c[14]), .y(y[14]));
  Leaf l15(.a(a[15]), .b(b[15]), .c(c[15]), .y(y[15]));
  Leaf l16(.a(a[16]), .b(b[16]), .c(c[16]), .y(y[16]));
  Leaf l17(.a(a[17]), .b(b[17]), .c(c[17]), .y(y[17]));
  Leaf l18(.a(a[18]), .b(b[18]), .c(c[18]), .y(y[18]));
  Leaf l19(.a(a[19]), .b(b[19]), .c(c[19]), .y(y[19]));
  Leaf l20(.a(a[20]), .b(b[20]), .c(c[20]), .y(y[20]));
  Leaf l21(.a(a[21]), .b(b[21]), .c(c[21]), .y(y[21]));
  Leaf l22(.a(a[22]), .b(b[22]), .c(c[22]), .y(y[22]));
  Leaf l23(.a(a[23]), .b(b[23]), .c(c[23]), .y(y[23]));
  Leaf l24(.a(a[24]), .b(b[24]), .c(c[24]), .y(y[24]));
  Leaf l25(.a(a[25]), .b(b[25]), .c(c[25]), .y(y[25]));
  Leaf l26(.a(a[26]), .b(b[26]), .c(c[26]), .y(y[26]));
  Leaf l27(.a(a[27]), .b(b[27]), .c(c[27]), .y(y[27]));
  Leaf l28(.a(a[28]), .b(b[28]), .c(c[28]), .y(y[28]));
  Leaf l29(.a(a[29]), .b(b[29]), .c(c[29]), .y(y[29]));
  Leaf l30(.a(a[30]), .b(b[30]), .c(c[30]), .y(y[30]));
  Leaf l31(.a(a[31]), .b(b[31]), .c(c[31]), .y(y[31]));
  Leaf l32(.a(a[32]), .b(b[32]), .c(c[32]), .y(y[32]));
  Leaf l33(.a(a[33]), .b(b[33]), .c(c[33]), .y(y[33]));
  Leaf l34(.a(a[34]), .b(b[34]), .c(c[34]), .y(y[34]));
  Leaf l35(.a(a[35]), .b(b[35]), .c(c[35]), .y(y[35]));
  Leaf l36(.a(a[36]), .b(b[36]), .c(c[36]), .y(y[36]));
  Leaf l37(.a(a[37]), .b(b[37]), .c(c[37]), .y(y[37]));
  Leaf l38(.a(a[38]), .b(b[38]), .c(c[38]), .y(y[38]));
  Leaf l39(.a(a[39]), .b(b[39]), .c(c[39]), .y(y[39]));
  Leaf l40(.a(a[40]), .b(b[40]), .c(c[40]), .y(y[40]));
  Leaf l41(.a(a[41]), .b(b[41]), .c(c[41]), .y(y[41]));
  Leaf l42(.a(a[42]), .b(b[42]), .c(c[42]), .y(y[42]));
  Leaf l43(.a(a[43]), .b(b[43]), .c(c[43]), .y(y[43]));
  Leaf l44(.a(a[44]), .b(b[44]), .c(c[44]), .y(y[44]));
  Leaf l45(.a(a[45]), .b(b[45]), .c(c[45]), .y(y[45]));
  Leaf l46(.a(a[46]), .b(b[46]), .c(c[46]), .y(y[46]));
  Leaf l47(.a(a[47]), .b(b[47]), .c(c[47]), .y(y[47]));
  Leaf l48(.a(a[48]), .b(b[48]), .c(c[48]), .y(y[48]));
  Leaf l49(.a(a[49]), .b(b[49]), .c(c[49]), .y(y[49]));
  Leaf l50(.a(a[50]), .b(b[50]), .c(c[50]), .y(y[50]));
  Leaf l51(.a(a[51]), .b(b[51]), .c(c[51]), .y(y[51]));
  Leaf l52(.a(a[52]), .b(b[52]), .c(c[52]), .y(y[52]));
  Leaf l53(.a(a[53]), .b(b[53]), .c(c[53]), .y(y[53]));
  Leaf l54(.a(a[54]), .b(b[54]), .c(c[54]), .y(y[54]));
  Leaf l55(.a(a[55]), .b(b[55]), .c(c[55]), .y(y[55]));
  Leaf l56(.a(a[56]), .b(b[56]), .c(c[56]), .y(y[56]));
  Leaf l57(.a(a[57]), .b(b[57]), .c(c[57]), .y(y[57]));
  Leaf l58(.a(a[58]), .b(b[58]), .c(c[58]), .y(y[58]));
  Leaf l59(.a(a[59]), .b(b[59]), .c(c[59]), .y(y[59]));
  Leaf l60(.a(a[60]), .b(b[60]), .c(c[60]), .y(y[60]));
  Leaf l61(.a(a[61]), .b(b[61]), .c(c[61]), .y(y[61]));
  Leaf l62(.a(a[62]), .b(b[62]), .c(c[62]), .y(y[62]));
  Leaf l63(.a(a[63]), .b(b[63]), .c(c[63]), .y(y[63]));
  Leaf l64(.a(a[64]), .b(b[64]), .c(c[64]), .y(y[64]));
  Leaf l65(.a(a[65]), .b(b[65]), .c(c[65]), .y(y[65]));
  Leaf l66(.a(a[66]), .b(b[66]), .c(c[66]), .y(y[66]));
  Leaf l67(.a(a[67]), .b(b[67]), .c(c[67]), .y(y[67]));
  Leaf l68(.a(a[68]), .b(b[68]), .c(c[68]), .y(y[68]));
  Leaf l69(.a(a[69]), .b(b[69]), .c(c[69]), .y(y[69]));
  Leaf l70(.a(a[70]), .b(b[70]), .c(c[70]), .y(y[70]));
  Leaf l71(.a(a[71]), .b(b[71]), .c(c[71]), .y(y[71]));
  Leaf l72(.a(a[72]), .b(b[72]), .c(c[72]), .y(y[72]));
  Leaf l73(.a(a[73]), .b(b[73]), .c(c[73]), .y(y[73]));
  Leaf l74(.a(a[74]), .b(b[74]), .c(c[74]), .y(y[74]));
  Leaf l75(.a(a[75]), .b(b[75]), .c(c[75]), .y(y[75]));
  Leaf l76(.a(a[76]), .b(b[76]), .c(c[76]), .y(y[76]));
  Leaf l77(.a(a[77]), .b(b[77]), .c(c[77]), .y(y[77]));
  Leaf l78(.a(a[78]), .b(b[78]), .c(c[78]), .y(y[78]));
  Leaf l79(.a(a[79]), .b(b[79]), .c(c[79]), .y(y[79]));
  Leaf l80(.a(a[80]), .b(b[80]), .c(c[80]), .y(y[80]));
  Leaf l81(.a(a[81]), .b(b[81]), .c(c[81]), .y(y[81]));
  Leaf l82(.a(a[82]), .b(b[82]), .c(c[82]), .y(y[82]));
  Leaf l83(.a(a[83]), .b(b[83]), .c(c[83]), .y(y[83]));
  Leaf l84(.a(a[84]), .b(b[84]), .c(c[84]), .y(y[84]));
  Leaf l85(.a(a[85]), .b(b[85]), .c(c[85]), .y(y[85]));
  Leaf l86(.a(a[86]), .b(b[86]), .c(c[86]), .y(y[86]));
  Leaf l87(.a(a[87]), .b(b[87]), .c(c[87]), .y(y[87]));
  Leaf l88(.a(a[88]), .b(b[88]), .c(c[88]), .y(y[88]));
  Leaf l89(.a(a[89]), .b(b[89]), .c(c[89]), .y(y[89]));
  Leaf l90(.a(a[90]), .b(b[90]), .c(c[90]), .y(y[90]));
  Leaf l91(.a(a[91]), .b(b[91]), .c(c[91]), .y(y[91]));
  Leaf l92(.a(a[92]), .b(b[92]), .c(c[92]), .y(y[92]));
  Leaf l93(.a(a[93]), .b(b[93]), .c(c[93]), .y(y[93]));
  Leaf l94(.a(a[94]), .b(b[94]), .c(c[94]), .y(y[94]));
  Leaf l95(.a(a[95]), .b(b[95]), .c(c[95]), .y(y[95]));
  Leaf l96(.a(a[96]), .b(b[96]), .c(c[96]), .y(y[96]));
  Leaf l97(.a(a[97]), .b(b[97]), .c(c[97]), .y(y[97]));
  Leaf l98(.a(a[98]), .b(b[98]), .c(c[98]), .y(y[98]));
  Leaf l99(.a(a[99]), .b(b[99]), .c(c[99]), .y(y[99]));
  Leaf l100(.a(a[100]), .b(b[100]), .c(c[100]), .y(y[100]));
  Leaf l101(.a(a[101]), .b(b[101]), .c(c[101]), .y(y[101]));
  Leaf l102(.a(a[102]), .b(b[102]), .c(c[102]), .y(y[102]));
  Leaf l103(.a(a[103]), .b(b[103]), .c(c[103]), .y(y[103]));
  Leaf l104(.a(a[104]), .b(b[104]), .c(c[104]), .y(y[104]));
  Leaf l105(.a(a[105]), .b(b[105]), .c(c[105]), .y(y[105]));
  Leaf l106(.a(a[106]), .b(b[106]), .c(c[106]), .y(y[106]));
  Leaf l107(.a(a[107]), .b(b[107]), .c(c[107]), .y(y[107]));
  Leaf l108(.a(a[108]), .b(b[108]), .c(c[108]), .y(y[108]));
  Leaf l109(.a(a[109]), .b(b[109]), .c(c[109]), .y(y[109]));
  Leaf l110(.a(a[110]), .b(b[110]), .c(c[110]), .y(y[110]));
  Leaf l111(.a(a[111]), .b(b[111]), .c(c[111]), .y(y[111]));
  Leaf l112(.a(a[112]), .b(b[112]), .c(c[112]), .y(y[112]));
  Leaf l113(.a(a[113]), .b(b[113]), .c(c[113]), .y(y[113]));
  Leaf l114(.a(a[114]), .b(b[114]), .c(c[114]), .y(y[114]));
  Leaf l115(.a(a[115]), .b(b[115]), .c(c[115]), .y(y[115]));
  Leaf l116(.a(a[116]), .b(b[116]), .c(c[116]), .y(y[116]));
  Leaf l117(.a(a[117]), .b(b[117]), .c(c[117]), .y(y[117]));
  Leaf l118(.a(a[118]), .b(b[118]), .c(c[118]), .y(y[118]));
  Leaf l119(.a(a[119]), .b(b[119]), .c(c[119]), .y(y[119]));
  Leaf l120(.a(a[120]), .b(b[120]), .c(c[120]), .y(y[120]));
  Leaf l121(.a(a[121]), .b(b[121]), .c(c[121]), .y(y[121]));
  Leaf l122(.a(a[122]), .b(b[122]), .c(c[122]), .y(y[122]));
  Leaf l123(.a(a[123]), .b(b[123]), .c(c[123]), .y(y[123]));
  Leaf l124(.a(a[124]), .b(b[124]), .c(c[124]), .y(y[124]));
  Leaf l125(.a(a[125]), .b(b[125]), .c(c[125]), .y(y[125]));
  Leaf l126(.a(a[126]), .b(b[126]), .c(c[126]), .y(y[126]));
  Leaf l127(.a(a[127]), .b(b[127]), .c(c[127]), .y(y[127]));
  Leaf l128(.a(a[128]), .b(b[128]), .c(c[128]), .y(y[128]));
  Leaf l129(.a(a[129]), .b(b[129]), .c(c[129]), .y(y[129]));
  Leaf l130(.a(a[130]), .b(b[130]), .c(c[130]), .y(y[130]));
  Leaf l131(.a(a[131]), .b(b[131]), .c(c[131]), .y(y[131]));
  Leaf l132(.a(a[132]), .b(b[132]), .c(c[132]), .y(y[132]));
  Leaf l133(.a(a[133]), .b(b[133]), .c(c[133]), .y(y[133]));
  Leaf l134(.a(a[134]), .b(b[134]), .c(c[134]), .y(y[134]));
  Leaf l135(.a(a[135]), .b(b[135]), .c(c[135]), .y(y[135]));
  Leaf l136(.a(a[136]), .b(b[136]), .c(c[136]), .y(y[136]));
  Leaf l137(.a(a[137]), .b(b[137]), .c(c[137]), .y(y[137]));
  Leaf l138(.a(a[138]), .b(b[138]), .c(c[138]), .y(y[138]));
  Leaf l139(.a(a[139]), .b(b[139]), .c(c[139]), .y(y[139]));
  Leaf l140(.a(a[140]), .b(b[140]), .c(c[140]), .y(y[140]));
  Leaf l141(.a(a[141]), .b(b[141]), .c(c[141]), .y(y[141]));
  Leaf l142(.a(a[142]), .b(b[142]), .c(c[142]), .y(y[142]));
  Leaf l143(.a(a[143]), .b(b[143]), .c(c[143]), .y(y[143]));
  Leaf l144(.a(a[144]), .b(b[144]), .c(c[144]), .y(y[144]));
  Leaf l145(.a(a[145]), .b(b[145]), .c(c[145]), .y(y[145]));
  Leaf l146(.a(a[146]), .b(b[146]), .c(c[146]), .y(y[146]));
  Leaf l147(.a(a[147]), .b(b[147]), .c(c[147]), .y(y[147]));
  Leaf l148(.a(a[148]), .b(b[148]), .c(c[148]), .y(y[148]));
  Leaf l149(.a(a[149]), .b(b[149]), .c(c[149]), .y(y[149]));
  Leaf l150(.a(a[150]), .b(b[150]), .c(c[150]), .y(y[150]));
  Leaf l151(.a(a[151]), .b(b[151]), .c(c[151]), .y(y[151]));
  Leaf l152(.a(a[152]), .b(b[152]), .c(c[152]), .y(y[152]));
  Leaf l153(.a(a[153]), .b(b[153]), .c(c[153]), .y(y[153]));
  Leaf l154(.a(a[154]), .b(b[154]), .c(c[154]), .y(y[154]));
  Leaf l155(.a(a[155]), .b(b[155]), .c(c[155]), .y(y[155]));
  Leaf l156(.a(a[156]), .b(b[156]), .c(c[156]), .y(y[156]));
  Leaf l157(.a(a[157]), .b(b[157]), .c(c[157]), .y(y[157]));
  Leaf l158(.a(a[158]), .b(b[158]), .c(c[158]), .y(y[158]));
  Leaf l159(.a(a[159]), .b(b[159]), .c(c[159]), .y(y[159]));
  Leaf l160(.a(a[160]), .b(b[160]), .c(c[160]), .y(y[160]));
  Leaf l161(.a(a[161]), .b(b[161]), .c(c[161]), .y(y[161]));
  Leaf l162(.a(a[162]), .b(b[162]), .c(c[162]), .y(y[162]));
  Leaf l163(.a(a[163]), .b(b[163]), .c(c[163]), .y(y[163]));
  Leaf l164(.a(a[164]), .b(b[164]), .c(c[164]), .y(y[164]));
  Leaf l165(.a(a[165]), .b(b[165]), .c(c[165]), .y(y[165]));
  Leaf l166(.a(a[166]), .b(b[166]), .c(c[166]), .y(y[166]));
  Leaf l167(.a(a[167]), .b(b[167]), .c(c[167]), .y(y[167]));
  Leaf l168(.a(a[168]), .b(b[168]), .c(c[168]), .y(y[168]));
  Leaf l169(.a(a[169]), .b(b[169]), .c(c[169]), .y(y[169]));
  Leaf l170(.a(a[170]), .b(b[170]), .c(c[170]), .y(y[170]));
  Leaf l171(.a(a[171]), .b(b[171]), .c(c[171]), .y(y[171]));
  Leaf l172(.a(a[172]), .b(b[172]), .c(c[172]), .y(y[172]));
  Leaf l173(.a(a[173]), .b(b[173]), .c(c[173]), .y(y[173]));
  Leaf l174(.a(a[174]), .b(b[174]), .c(c[174]), .y(y[174]));
  Leaf l175(.a(a[175]), .b(b[175]), .c(c[175]), .y(y[175]));
  Leaf l176(.a(a[176]), .b(b[176]), .c(c[176]), .y(y[176]));
  Leaf l177(.a(a[177]), .b(b[177]), .c(c[177]), .y(y[177]));
  Leaf l178(.a(a[178]), .b(b[178]), .c(c[178]), .y(y[178]));
  Leaf l179(.a(a[179]), .b(b[179]), .c(c[179]), .y(y[179]));
  Leaf l180(.a(a[180]), .b(b[180]), .c(c[180]), .y(y[180]));
  Leaf l181(.a(a[181]), .b(b[181]), .c(c[181]), .y(y[181]));
  Leaf l182(.a(a[182]), .b(b[182]), .c(c[182]), .y(y[182]));
  Leaf l183(.a(a[183]), .b(b[183]), .c(c[183]), .y(y[183]));
  Leaf l184(.a(a[184]), .b(b[184]), .c(c[184]), .y(y[184]));
  Leaf l185(.a(a[185]), .b(b[185]), .c(c[185]), .y(y[185]));
  Leaf l186(.a(a[186]), .b(b[186]), .c(c[186]), .y(y[186]));
  Leaf l187(.a(a[187]), .b(b[187]), .c(c[187]), .y(y[187]));
  Leaf l188(.a(a[188]), .b(b[188]), .c(c[188]), .y(y[188]));
  Leaf l189(.a(a[189]), .b(b[189]), .c(c[189]), .y(y[189]));
  Leaf l190(.a(a[190]), .b(b[190]), .c(c[190]), .y(y[190]));
  Leaf l191(.a(a[191]), .b(b[191]), .c(c[191]), .y(y[191]));
  Leaf l192(.a(a[192]), .b(b[192]), .c(c[192]), .y(y[192]));
  Leaf l193(.a(a[193]), .b(b[193]), .c(c[193]), .y(y[193]));
  Leaf l194(.a(a[194]), .b(b[194]), .c(c[194]), .y(y[194]));
  Leaf l195(.a(a[195]), .b(b[195]), .c(c[195]), .y(y[195]));
  Leaf l196(.a(a[196]), .b(b[196]), .c(c[196]), .y(y[196]));
  Leaf l197(.a(a[197]), .b(b[197]), .c(c[197]), .y(y[197]));
  Leaf l198(.a(a[198]), .b(b[198]), .c(c[198]), .y(y[198]));
  Leaf l199(.a(a[199]), .b(b[199]), .c(c[199]), .y(y[199]));
  Leaf l200(.a(a[200]), .b(b[200]), .c(c[200]), .y(y[200]));
  Leaf l201(.a(a[201]), .b(b[201]), .c(c[201]), .y(y[201]));
  Leaf l202(.a(a[202]), .b(b[202]), .c(c[202]), .y(y[202]));
  Leaf l203(.a(a[203]), .b(b[203]), .c(c[203]), .y(y[203]));
  Leaf l204(.a(a[204]), .b(b[204]), .c(c[204]), .y(y[204]));
  Leaf l205(.a(a[205]), .b(b[205]), .c(c[205]), .y(y[205]));
  Leaf l206(.a(a[206]), .b(b[206]), .c(c[206]), .y(y[206]));
  Leaf l207(.a(a[207]), .b(b[207]), .c(c[207]), .y(y[207]));
  Leaf l208(.a(a[208]), .b(b[208]), .c(c[208]), .y(y[208]));
  Leaf l209(.a(a[209]), .b(b[209]), .c(c[209]), .y(y[209]));
  Leaf l210(.a(a[210]), .b(b[210]), .c(c[210]), .y(y[210]));
  Leaf l211(.a(a[211]), .b(b[211]), .c(c[211]), .y(y[211]));
  Leaf l212(.a(a[212]), .b(b[212]), .c(c[212]), .y(y[212]));
  Leaf l213(.a(a[213]), .b(b[213]), .c(c[213]), .y(y[213]));
  Leaf l214(.a(a[214]), .b(b[214]), .c(c[214]), .y(y[214]));
  Leaf l215(.a(a[215]), .b(b[215]), .c(c[215]), .y(y[215]));
  Leaf l216(.a(a[216]), .b(b[216]), .c(c[216]), .y(y[216]));
  Leaf l217(.a(a[217]), .b(b[217]), .c(c[217]), .y(y[217]));
  Leaf l218(.a(a[218]), .b(b[218]), .c(c[218]), .y(y[218]));
  Leaf l219(.a(a[219]), .b(b[219]), .c(c[219]), .y(y[219]));
  Leaf l220(.a(a[220]), .b(b[220]), .c(c[220]), .y(y[220]));
  Leaf l221(.a(a[221]), .b(b[221]), .c(c[221]), .y(y[221]));
  Leaf l222(.a(a[222]), .b(b[222]), .c(c[222]), .y(y[222]));
  Leaf l223(.a(a[223]), .b(b[223]), .c(c[223]), .y(y[223]));
  Leaf l224(.a(a[224]), .b(b[224]), .c(c[224]), .y(y[224]));
  Leaf l225(.a(a[225]), .b(b[225]), .c(c[225]), .y(y[225]));
  Leaf l226(.a(a[226]), .b(b[226]), .c(c[226]), .y(y[226]));
  Leaf l227(.a(a[227]), .b(b[227]), .c(c[227]), .y(y[227]));
  Leaf l228(.a(a[228]), .b(b[228]), .c(c[228]), .y(y[228]));
  Leaf l229(.a(a[229]), .b(b[229]), .c(c[229]), .y(y[229]));
  Leaf l230(.a(a[230]), .b(b[230]), .c(c[230]), .y(y[230]));
  Leaf l231(.a(a[231]), .b(b[231]), .c(c[231]), .y(y[231]));
  Leaf l232(.a(a[232]), .b(b[232]), .c(c[232]), .y(y[232]));
  Leaf l233(.a(a[233]), .b(b[233]), .c(c[233]), .y(y[233]));
  Leaf l234(.a(a[234]), .b(b[234]), .c(c[234]), .y(y[234]));
  Leaf l235(.a(a[235]), .b(b[235]), .c(c[235]), .y(y[235]));
  Leaf l236(.a(a[236]), .b(b[236]), .c(c[236]), .y(y[236]));
  Leaf l237(.a(a[237]), .b(b[237]), .c(c[237]), .y(y[237]));
  Leaf l238(.a(a[238]), .b(b[238]), .c(c[238]), .y(y[238]));
  Leaf l239(.a(a[239]), .b(b[239]), .c(c[239]), .y(y[239]));
  Leaf l240(.a(a[240]), .b(b[240]), .c(c[240]), .y(y[240]));
  Leaf l241(.a(a[241]), .b(b[241]), .c(c[241]), .y(y[241]));
  Leaf l242(.a(a[242]), .b(b[242]), .c(c[242]), .y(y[242]));
  Leaf l243(.a(a[243]), .b(b[243]), .c(c[243]), .y(y[243]));
  Leaf l244(.a(a[244]), .b(b[244]), .c(c[244]), .y(y[244]));
  Leaf l245(.a(a[245]), .b(b[245]), .c(c[245]), .y(y[245]));
  Leaf l246(.a(a[246]), .b(b[246]), .c(c[246]), .y(y[246]));
  Leaf l247(.a(a[247]), .b(b[247]), .c(c[247]), .y(y[247]));
  Leaf l248(.a(a[248]), .b(b[248]), .c(c[248]), .y(y[248]));
  Leaf l249(.a(a[249]), .b(b[249]), .c(c[249]), .y(y[249]));
  Leaf l250(.a(a[250]), .b(b[250]), .c(c[250]), .y(y[250]));
  Leaf l251(.a(a[251]), .b(b[251]), .c(c[251]), .y(y[251]));
  Leaf l252(.a(a[252]), .b(b[252]), .c(c[252]), .y(y[252]));
  Leaf l253(.a(a[253]), .b(b[253]), .c(c[253]), .y(y[253]));
  Leaf l254(.a(a[254]), .b(b[254]), .c(c[254]), .y(y[254]));
  Leaf l255(.a(a[255]), .b(b[255]), .c(c[255]), .y(y[255]));
endmodule

module TopLarge(input [16383:0] a, input [16383:0] b, input [16383:0] c, output [16383:0] y);
  Mid m0(.a(a[255:0]), .b(b[255:0]), .c(c[255:0]), .y(y[255:0]));
  Mid m1(.a(a[511:256]), .b(b[511:256]), .c(c[511:256]), .y(y[511:256]));
  Mid m2(.a(a[767:512]), .b(b[767:512]), .c(c[767:512]), .y(y[767:512]));
  Mid m3(.a(a[1023:768]), .b(b[1023:768]), .c(c[1023:768]), .y(y[1023:768]));
  Mid m4(.a(a[1279:1024]), .b(b[1279:1024]), .c(c[1279:1024]), .y(y[1279:1024]));
  Mid m5(.a(a[1535:1280]), .b(b[1535:1280]), .c(c[1535:1280]), .y(y[1535:1280]));
  Mid m6(.a(a[1791:1536]), .b(b[1791:1536]), .c(c[1791:1536]), .y(y[1791:1536]));
  Mid m7(.a(a[2047:1792]), .b(b[2047:1792]), .c(c[2047:1792]), .y(y[2047:1792]));
  Mid m8(.a(a[2303:2048]), .b(b[2303:2048]), .c(c[2303:2048]), .y(y[2303:2048]));
  Mid m9(.a(a[2559:2304]), .b(b[2559:2304]), .c(c[2559:2304]), .y(y[2559:2304]));
  Mid m10(.a(a[2815:2560]), .b(b[2815:2560]), .c(c[2815:2560]), .y(y[2815:2560]));
  Mid m11(.a(a[3071:2816]), .b(b[3071:2816]), .c(c[3071:2816]), .y(y[3071:2816]));
  Mid m12(.a(a[3327:3072]), .b(b[3327:3072]), .c(c[3327:3072]), .y(y[3327:3072]));
  Mid m13(.a(a[3583:3328]), .b(b[3583:3328]), .c(c[3583:3328]), .y(y[3583:3328]));
  Mid m14(.a(a[3839:3584]), .b(b[3839:3584]), .c(c[3839:3584]), .y(y[3839:3584]));
  Mid m15(.a(a[4095:3840]), .b(b[4095:3840]), .c(c[4095:3840]), .y(y[4095:3840]));
  Mid m16(.a(a[4351:4096]), .b(b[4351:4096]), .c(c[4351:4096]), .y(y[4351:4096]));
  Mid m17(.a(a[4607:4352]), .b(b[4607:4352]), .c(c[4607:4352]), .y(y[4607:4352]));
  Mid m18(.a(a[4863:4608]), .b(b[4863:4608]), .c(c[4863:4608]), .y(y[4863:4608]));
  Mid m19(.a(a[5119:4864]), .b(b[5119:4864]), .c(c[5119:4864]), .y(y[5119:4864]));
  Mid m20(.a(a[5375:5120]), .b(b[5375:5120]), .c(c[5375:5120]), .y(y[5375:5120]));
  Mid m21(.a(a[5631:5376]), .b(b[5631:5376]), .c(c[5631:5376]), .y(y[5631:5376]));
  Mid m22(.a(a[5887:5632]), .b(b[5887:5632]), .c(c[5887:5632]), .y(y[5887:5632]));
  Mid m23(.a(a[6143:5888]), .b(b[6143:5888]), .c(c[6143:5888]), .y(y[6143:5888]));
  Mid m24(.a(a[6399:6144]), .b(b[6399:6144]), .c(c[6399:6144]), .y(y[6399:6144]));
  Mid m25(.a(a[6655:6400]), .b(b[6655:6400]), .c(c[6655:6400]), .y(y[6655:6400]));
  Mid m26(.a(a[6911:6656]), .b(b[6911:6656]), .c(c[6911:6656]), .y(y[6911:6656]));
  Mid m27(.a(a[7167:6912]), .b(b[7167:6912]), .c(c[7167:6912]), .y(y[7167:6912]));
  Mid m28(.a(a[7423:7168]), .b(b[7423:7168]), .c(c[7423:7168]), .y(y[7423:7168]));
  Mid m29(.a(a[7679:7424]), .b(b[7679:7424]), .c(c[7679:7424]), .y(y[7679:7424]));
  Mid m30(.a(a[7935:7680]), .b(b[7935:7680]), .c(c[7935:7680]), .y(y[7935:7680]));
  Mid m31(.a(a[8191:7936]), .b(b[8191:7936]), .c(c[8191:7936]), .y(y[8191:7936]));
  Mid m32(.a(a[8447:8192]), .b(b[8447:8192]), .c(c[8447:8192]), .y(y[8447:8192]));
  Mid m33(.a(a[8703:8448]), .b(b[8703:8448]), .c(c[8703:8448]), .y(y[8703:8448]));
  Mid m34(.a(a[8959:8704]), .b(b[8959:8704]), .c(c[8959:8704]), .y(y[8959:8704]));
  Mid m35(.a(a[9215:8960]), .b(b[9215:8960]), .c(c[9215:8960]), .y(y[9215:8960]));
  Mid m36(.a(a[9471:9216]), .b(b[9471:9216]), .c(c[9471:9216]), .y(y[9471:9216]));
  Mid m37(.a(a[9727:9472]), .b(b[9727:9472]), .c(c[9727:9472]), .y(y[9727:9472]));
  Mid m38(.a(a[9983:9728]), .b(b[9983:9728]), .c(c[9983:9728]), .y(y[9983:9728]));
  Mid m39(.a(a[10239:9984]), .b(b[10239:9984]), .c(c[10239:9984]), .y(y[10239:9984]));
  Mid m40(.a(a[10495:10240]), .b(b[10495:10240]), .c(c[10495:10240]), .y(y[10495:10240]));
  Mid m41(.a(a[10751:10496]), .b(b[10751:10496]), .c(c[10751:10496]), .y(y[10751:10496]));
  Mid m42(.a(a[11007:10752]), .b(b[11007:10752]), .c(c[11007:10752]), .y(y[11007:10752]));
  Mid m43(.a(a[11263:11008]), .b(b[11263:11008]), .c(c[11263:11008]), .y(y[11263:11008]));
  Mid m44(.a(a[11519:11264]), .b(b[11519:11264]), .c(c[11519:11264]), .y(y[11519:11264]));
  Mid m45(.a(a[11775:11520]), .b(b[11775:11520]), .c(c[11775:11520]), .y(y[11775:11520]));
  Mid m46(.a(a[12031:11776]), .b(b[12031:11776]), .c(c[12031:11776]), .y(y[12031:11776]));
  Mid m47(.a(a[12287:12032]), .b(b[12287:12032]), .c(c[12287:12032]), .y(y[12287:12032]));
  Mid m48(.a(a[12543:12288]), .b(b[12543:12288]), .c(c[12543:12288]), .y(y[12543:12288]));
  Mid m49(.a(a[12799:12544]), .b(b[12799:12544]), .c(c[12799:12544]), .y(y[12799:12544]));
  Mid m50(.a(a[13055:12800]), .b(b[13055:12800]), .c(c[13055:12800]), .y(y[13055:12800]));
  Mid m51(.a(a[13311:13056]), .b(b[13311:13056]), .c(c[13311:13056]), .y(y[13311:13056]));
  Mid m52(.a(a[13567:13312]), .b(b[13567:13312]), .c(c[13567:13312]), .y(y[13567:13312]));
  Mid m53(.a(a[13823:13568]), .b(b[13823:13568]), .c(c[13823:13568]), .y(y[13823:13568]));
  Mid m54(.a(a[14079:13824]), .b(b[14079:13824]), .c(c[14079:13824]), .y(y[14079:13824]));
  Mid m55(.a(a[14335:14080]), .b(b[14335:14080]), .c(c[14335:14080]), .y(y[14335:14080]));
  Mid m56(.a(a[14591:14336]), .b(b[14591:14336]), .c(c[14591:14336]), .y(y[14591:14336]));
  Mid m57(.a(a[14847:14592]), .b(b[14847:14592]), .c(c[14847:14592]), .y(y[14847:14592]));
  Mid m58(.a(a[15103:14848]), .b(b[15103:14848]), .c(c[15103:14848]), .y(y[15103:14848]));
  Mid m59(.a(a[15359:15104]), .b(b[15359:15104]), .c(c[15359:15104]), .y(y[15359:15104]));
  Mid m60(.a(a[15615:15360]), .b(b[15615:15360]), .c(c[15615:15360]), .y(y[15615:15360]));
  Mid m61(.a(a[15871:15616]), .b(b[15871:15616]), .c(c[15871:15616]), .y(y[15871:15616]));
  Mid m62(.a(a[16127:15872]), .b(b[16127:15872]), .c(c[16127:15872]), .y(y[16127:15872]));
  Mid m63(.a(a[16383:16128]), .b(b[16383:16128]), .c(c[16383:16128]), .y(y[16383:16128]));
endmodule
