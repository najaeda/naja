// SPDX-FileCopyrightText: 2026 The Naja authors <https://github.com/najaeda/naja/blob/main/AUTHORS>
//
// SPDX-License-Identifier: Apache-2.0

module byte_ports_top(
  input byte a,
  output byte y
);
  assign y = a;
endmodule
