module \#model0 (input \%t0 , input \12t1@ , input [3:0] \3 4 , input [-5:2] \## );
endmodule //#model0

module \design@ ();
\#model0  \0ins  (
  .\%t0 (),
  .\12t1@ (),
  .\3 4 (),
  .\## ()
);
endmodule //design@
