// SPDX-FileCopyrightText: 2026 The Naja authors <https://github.com/najaeda/naja/blob/main/AUTHORS>
//
// SPDX-License-Identifier: Apache-2.0

module implicit_width_ports_top(
  input int wide_i,
  input bit bit_i,
  output int wide_o
);
endmodule
