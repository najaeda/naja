////////////////////////////////////////////////////////////////////////////////
#IGNORE#
#IGNORE#
#IGNORE#
#IGNORE#
////////////////////////////////////////////////////////////////////////////////

module top_bus_assign_compression();
wire [3:0] source_bus;
wire [3:0] sink_bus;

assign sink_bus = source_bus;
endmodule //top_bus_assign_compression
