// SPDX-FileCopyrightText: 2026 The Naja authors <https://github.com/najaeda/naja/blob/main/AUTHORS>
//
// SPDX-License-Identifier: Apache-2.0

module compatible_net_scalar_mismatch_top(
  input logic a,
  input logic b,
  output logic y
);
  logic [1:0] and_y;
  assign y = a & b;
endmodule
