/*
  Testing empty connection
*/

module test_empty_instance_connection();
  model0 inst0(.A());
endmodule