module seq_list_single_empty_stmt_unsupported(
  input logic clk,
  output logic q
);
  // Single-item statement list with an empty statement.
  always begin
    ;
  end
endmodule
